* File: inv.pex.netlist.sp
* Created: Wed Oct 20 00:03:58 2021
* Program "Calibre xRC"
* Version "v2012.2_36.25"
* 
*----------------------------------------------------------------------
* Paramters and models 
*----------------------------------------------------------------------
.param SUPPLY=3.3
.include "tsmc_018_pex.sp"
.temp 70
.option post
*----------------------------------------------------------------------
.include "inv.pex.netlist"
*----------------------------------------------------------------------
* Simulation netlist 
*----------------------------------------------------------------------
Vdd  vdd  gnd 'SUPPLY'
Vin vin gnd PULSE 0 'SUPPLY' 25ps 0ps 0ps 35ps 80ps
X1 vin vout gnd vdd INV
*----------------------------------------------------------------------
* Stimulus 
*----------------------------------------------------------------------
.tran 0.1ps 80ps
.end
*